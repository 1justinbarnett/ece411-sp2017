package lc3b_config;

parameter USE_ADVANCED_CACHE = 1;
parameter USE_VICTIM_CACHES = 1;
parameter USE_BRANCH_PREDICTION = 1;

endpackage : lc3b_config
